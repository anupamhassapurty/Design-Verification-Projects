library verilog;
use verilog.vl_types.all;
entity lod_test is
end lod_test;

library verilog;
use verilog.vl_types.all;
entity muxa is
    port(
        s               : in     vl_logic;
        y               : out    vl_logic
    );
end muxa;
